// rippleUpTop.v

`include "rippleUp.v"

module testBench;

endmodule

module Tester();

endmodule