library verilog;
use verilog.vl_types.all;
entity DownCounterSchematic_vlg_vec_tst is
end DownCounterSchematic_vlg_vec_tst;
