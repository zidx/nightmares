library verilog;
use verilog.vl_types.all;
entity DownCounterSchematic_vlg_check_tst is
    port(
        PIN_V16         : in     vl_logic;
        PIN_V17         : in     vl_logic;
        PIN_V18         : in     vl_logic;
        PIN_W16         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end DownCounterSchematic_vlg_check_tst;
