library verilog;
use verilog.vl_types.all;
entity DE1_SoC is
    generic(
        blank           : vl_logic_vector(0 to 6) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        fiveSec         : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        sevenSec        : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        eightSec        : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        whichClock      : integer := 6
    );
    port(
        CLOCK_50        : in     vl_logic;
        HEX0            : out    vl_logic_vector(6 downto 0);
        HEX1            : out    vl_logic_vector(6 downto 0);
        HEX2            : out    vl_logic_vector(6 downto 0);
        HEX3            : out    vl_logic_vector(6 downto 0);
        HEX4            : out    vl_logic_vector(6 downto 0);
        HEX5            : out    vl_logic_vector(6 downto 0);
        KEY             : in     vl_logic_vector(3 downto 0);
        LEDR            : out    vl_logic_vector(9 downto 0);
        SW              : in     vl_logic_vector(9 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of blank : constant is 1;
    attribute mti_svvh_generic_type of fiveSec : constant is 1;
    attribute mti_svvh_generic_type of sevenSec : constant is 1;
    attribute mti_svvh_generic_type of eightSec : constant is 1;
    attribute mti_svvh_generic_type of whichClock : constant is 1;
end DE1_SoC;
