library verilog;
use verilog.vl_types.all;
entity switchesqsys_mm_interconnect_0_cmd_demux_001 is
    port(
        sink_valid      : in     vl_logic_vector(0 downto 0);
        sink_data       : in     vl_logic_vector(91 downto 0);
        sink_channel    : in     vl_logic_vector(11 downto 0);
        sink_startofpacket: in     vl_logic;
        sink_endofpacket: in     vl_logic;
        sink_ready      : out    vl_logic;
        src0_valid      : out    vl_logic;
        src0_data       : out    vl_logic_vector(91 downto 0);
        src0_channel    : out    vl_logic_vector(11 downto 0);
        src0_startofpacket: out    vl_logic;
        src0_endofpacket: out    vl_logic;
        src0_ready      : in     vl_logic;
        src1_valid      : out    vl_logic;
        src1_data       : out    vl_logic_vector(91 downto 0);
        src1_channel    : out    vl_logic_vector(11 downto 0);
        src1_startofpacket: out    vl_logic;
        src1_endofpacket: out    vl_logic;
        src1_ready      : in     vl_logic;
        src2_valid      : out    vl_logic;
        src2_data       : out    vl_logic_vector(91 downto 0);
        src2_channel    : out    vl_logic_vector(11 downto 0);
        src2_startofpacket: out    vl_logic;
        src2_endofpacket: out    vl_logic;
        src2_ready      : in     vl_logic;
        src3_valid      : out    vl_logic;
        src3_data       : out    vl_logic_vector(91 downto 0);
        src3_channel    : out    vl_logic_vector(11 downto 0);
        src3_startofpacket: out    vl_logic;
        src3_endofpacket: out    vl_logic;
        src3_ready      : in     vl_logic;
        src4_valid      : out    vl_logic;
        src4_data       : out    vl_logic_vector(91 downto 0);
        src4_channel    : out    vl_logic_vector(11 downto 0);
        src4_startofpacket: out    vl_logic;
        src4_endofpacket: out    vl_logic;
        src4_ready      : in     vl_logic;
        src5_valid      : out    vl_logic;
        src5_data       : out    vl_logic_vector(91 downto 0);
        src5_channel    : out    vl_logic_vector(11 downto 0);
        src5_startofpacket: out    vl_logic;
        src5_endofpacket: out    vl_logic;
        src5_ready      : in     vl_logic;
        src6_valid      : out    vl_logic;
        src6_data       : out    vl_logic_vector(91 downto 0);
        src6_channel    : out    vl_logic_vector(11 downto 0);
        src6_startofpacket: out    vl_logic;
        src6_endofpacket: out    vl_logic;
        src6_ready      : in     vl_logic;
        src7_valid      : out    vl_logic;
        src7_data       : out    vl_logic_vector(91 downto 0);
        src7_channel    : out    vl_logic_vector(11 downto 0);
        src7_startofpacket: out    vl_logic;
        src7_endofpacket: out    vl_logic;
        src7_ready      : in     vl_logic;
        src8_valid      : out    vl_logic;
        src8_data       : out    vl_logic_vector(91 downto 0);
        src8_channel    : out    vl_logic_vector(11 downto 0);
        src8_startofpacket: out    vl_logic;
        src8_endofpacket: out    vl_logic;
        src8_ready      : in     vl_logic;
        src9_valid      : out    vl_logic;
        src9_data       : out    vl_logic_vector(91 downto 0);
        src9_channel    : out    vl_logic_vector(11 downto 0);
        src9_startofpacket: out    vl_logic;
        src9_endofpacket: out    vl_logic;
        src9_ready      : in     vl_logic;
        src10_valid     : out    vl_logic;
        src10_data      : out    vl_logic_vector(91 downto 0);
        src10_channel   : out    vl_logic_vector(11 downto 0);
        src10_startofpacket: out    vl_logic;
        src10_endofpacket: out    vl_logic;
        src10_ready     : in     vl_logic;
        src11_valid     : out    vl_logic;
        src11_data      : out    vl_logic_vector(91 downto 0);
        src11_channel   : out    vl_logic_vector(11 downto 0);
        src11_startofpacket: out    vl_logic;
        src11_endofpacket: out    vl_logic;
        src11_ready     : in     vl_logic;
        clk             : in     vl_logic;
        reset           : in     vl_logic
    );
end switchesqsys_mm_interconnect_0_cmd_demux_001;
